`include "def.v"
module LSB (
    input wire clk_in,
    input wire rst_in,
    input wire rdy_in,
    input wire clear,
    
    //REGFile
    
);
    
endmodule